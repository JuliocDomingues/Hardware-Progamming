library ieee;
use ieee.std_logic_1164.all;

entity tb_fulladder4 is
end;

architecture behavioral of tb_fulladder4 is
  signal 
